module libraw

import libs.libraw.c as _
