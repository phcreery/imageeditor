module common

// TODO rename to BackendID
pub enum DeviceMemoryContext {
	cpu
	cl
}
