module stb

// note, this will cause collision with vlang's stdlib stb module
#flag -I @VMODROOT/thirdparty/stb
