module write

#flag -I @VMODROOT/thirdparty/stb
#define STB_IMAGE_WRITE_IMPLEMENTATION
#include "stb_image_write.h"
