module main

pub fn print_console_header(version string) {
	println("
 ███████████  █████ ██████████
░░███░░░░░███░░███ ░░███░░░░░█
 ░███    ░███ ░███  ░███  █ ░ 
 ░██████████  ░███  ░██████   
 ░███░░░░░░   ░███  ░███░░█   
 ░███         ░███  ░███ ░   █
 █████        █████ ██████████
░░░░░        ░░░░░ ░░░░░░░░░░ 
                              
PEYTON'S IMAGE EDITOR v${version}
")
}
