module cimgui

import libs.cimgui.c as _
